-- This is your top level VHDL module

library IEEE;
use IEEE.std_logic_1164.all;

entity top is
  port(
    CLK   : in std_logic;
    RESET : in std_logic
  );
end entity top;

architecture Behavioral of top is
begin

end Behavioral;
